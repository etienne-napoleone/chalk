module chalk

const(
    Styles = {
        'bold': '1'
        'dim': '2'
        'underline': '4'
        'blink': '5'
        'reverse': '7'
        'hidden': '8'
    }
)
